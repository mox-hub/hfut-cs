library verilog;
use verilog.vl_types.all;
entity ram_tb is
end ram_tb;
