library verilog;
use verilog.vl_types.all;
entity alu_tb is
end alu_tb;
